module ARM(
    clk, rst
)


endmodule