library verilog;
use verilog.vl_types.all;
entity c17 is
    port(
        N1              : in     vl_logic;
        N2              : in     vl_logic;
        N3              : in     vl_logic;
        N6              : in     vl_logic;
        N7              : in     vl_logic;
        N22             : out    vl_logic;
        N23             : out    vl_logic
    );
end c17;
