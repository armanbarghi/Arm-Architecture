library verilog;
use verilog.vl_types.all;
entity ARM_TB is
end ARM_TB;
