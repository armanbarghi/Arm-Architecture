library verilog;
use verilog.vl_types.all;
entity Q_ARM_Testbench is
end Q_ARM_Testbench;
