library verilog;
use verilog.vl_types.all;
entity mytb is
end mytb;
