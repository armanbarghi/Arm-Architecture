library verilog;
use verilog.vl_types.all;
entity ARM_Testbench is
end ARM_Testbench;
