module IF_Stage_Reg(input clk, rst, freeze, flush,
                input [31:0] PC,
                output reg [31:0] PC, Inst);

endmodule
