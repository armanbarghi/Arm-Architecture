module InstMemory (
	AddrIn,
	Inst
);
	input [31:0] AddrIn;
	output [31:0] Inst;

	reg [31:0] mem[0:65535];

	initial begin
		// $readmemb("../Codes/InstMem.txt", mem);
		mem[0] = 32'b1110_00_1_1101_0_0000_0000_000000010100; //MOV R0 ,#20 //R0 = 20
		mem[1] = 32'b1110_00_1_1101_0_0000_0001_101000000001; //MOV R1 ,#4096 //R1 = 4096
		mem[2] = 32'b1110_00_1_1101_0_0000_0010_000100000011; //MOV R2 ,#0xC0000000 //R2 = -1073741824
		mem[3] = 32'b1110_00_0_0100_1_0010_0011_000000000010; //ADDS R3 ,R2,R2 //R3 = -2147483648 
		mem[4] = 32'b1110_00_0_0101_0_0000_0100_000000000000; //ADC R4 ,R0,R0 //R4 = 41
		mem[5] = 32'b1110_00_0_0010_0_0100_0101_000100000100; //SUB R5 ,R4,R4,LSL #2 //R5 = -123
		mem[6] = 32'b1110_00_0_0110_0_0000_0110_000010100000; //SBC R6 ,R0,R0,LSR #1 //R6 = 10
		mem[7] = 32'b1110_00_0_1100_0_0101_0111_000101000010; //ORR R7 ,R5,R2,ASR #2 //R7 = -123
		mem[8] = 32'b1110_00_0_0000_0_0111_1000_000000000011; //AND R8 ,R7,R3 //R8 = -2147483648
		mem[9] = 32'b1110_00_0_1111_0_0000_1001_000000000110; //MVN R9 ,R6 //R9 = -11
		mem[10] = 32'b1110_00_0_0001_0_0100_1010_000000000101; //EOR R10,R4,R5 //R10 = -84
		mem[11] = 32'b1110_00_0_1010_1_1000_0000_000000000110; //CMP R8 ,R6
		mem[12] = 32'b0001_00_0_0100_0_0001_0001_000000000001; //ADDNE R1 ,R1,R1 //R1 = 8192
		mem[13] = 32'b1110_00_0_1000_1_1001_0000_000000001000; //TST R9 ,R8
		mem[14] = 32'b0000_00_0_0100_0_0010_0010_000000000010; //ADDEQ R2 ,R2,R2 //R2 = -1073741824
		mem[15] = 32'b1110_00_1_1101_0_0000_0000_101100000001; //MOV R0 ,#1024 //R0 = 1024
		mem[16] = 32'b1110_01_0_0100_0_0000_0001_000000000000; //STR R1 ,[R0],#0 //MEM[1024] = 8192
     	mem[17] = 32'b1110_01_0_0100_1_0000_1011_000000000000; //LDR R11,[R0],#0 //R11 = 8192
     	mem[18] = 32'b1110_01_0_0100_0_0000_0010_000000000100; //STR R2 ,[R0],#4 //MEM[1028] = -1073741824
     	mem[19] = 32'b1110_01_0_0100_0_0000_0011_000000001000; //STR R3 ,[R0],#8 //MEM[1032] = -2147483648
     	mem[20] = 32'b1110_01_0_0100_0_0000_0100_000000001101; //STR R4 ,[R0],#13 //MEM[1036] = 41
     	mem[21] = 32'b1110_01_0_0100_0_0000_0101_000000010000; //STR R5 ,[R0],#16 //MEM[1040] = -123
     	mem[22] = 32'b1110_01_0_0100_0_0000_0110_000000010100; //STR R6 ,[R0],#20 //MEM[1044] = 10
     	mem[23] = 32'b1110_01_0_0100_1_0000_1010_000000000100; //LDR R10,[R0],#4 //R10 = -1073741824
     	mem[24] = 32'b1110_01_0_0100_0_0000_0111_000000011000; //STR R7 ,[R0],#24 //MEM[1048] = -123
     	mem[25] = 32'b1110_00_1_1101_0_0000_0001_000000000101; //MOV R1 ,#5 //R1 = 5
     	mem[26] = 32'b1110_00_1_1101_0_0000_0010_000000000000; //MOV R2 ,#0 //R2 = 0

     	// mem[27] = 32'b1110_00_1_1101_0_0000_0011_000000000000; //MOV R3 ,#0 //R3 = 0
     	// mem[28] = 32'b1110_00_0_0100_0_0000_0100_000100000011; //ADD R4 ,R0,R3,LSL #2
     	// mem[29] = 32'b1110_01_0_0100_1_0100_0101_000000000000; //LDR R5 ,[R4],#0
     	// mem[30] = 32'b1110_01_0_0100_1_0100_0110_000000000100; //LDR R6 ,[R4],#4
     	// mem[31] = 32'b1110_00_0_1010_1_0101_0000_000000000110; //CMP R5 ,R6
     	// mem[32] = 32'b1100_01_0_0100_0_0100_0110_000000000000; //STRGT R6 ,[R4],#0
     	// mem[33] = 32'b1100_01_0_0100_0_0100_0101_000000000100; //STRGT R5 ,[R4],#4
     	// mem[34] = 32'b1110_00_1_0100_0_0011_0011_000000000001; //ADD R3 ,R3,#1
		// mem[35] = 32'b1110_00_1_1010_1_0011_0000_000000000110; //CMP R3 ,#6
		// mem[36] = 32'b1011_10_1_0_111111111111111111110111 ;   //BLT #-9
		// mem[37] = 32'b1110_00_1_0100_0_0010_0010_000000000001; //ADD R2 ,R2,#1
		// mem[38] = 32'b1110_00_0_1010_1_0010_0000_000000000001; //CMP R2 ,R1
		// mem[39] = 32'b1011_10_1_0_111111111111111111110011 ;   //BLT #-13

		// mem[40] = 32'b1110_01_0_0100_1_0000_0001_000000000000; //LDR R1 ,[R0],#0 //R1 = -2147483648
		// mem[41] = 32'b1110_01_0_0100_1_0000_0010_000000000100; //LDR R2 ,[R0],#4 //R2 = -1073741824
		// mem[42] = 32'b1110_01_0_0100_1_0000_0011_000000001000; //LDR R3 ,[R0],#8 //R3 = -123
		// mem[43] = 32'b1110_01_0_0100_1_0000_0100_000000001100; //LDR R4 ,[R0],#12 //R4 = -123
		// mem[44] = 32'b1110_01_0_0100_1_0000_0101_000000010000; //LDR R5 ,[R0],#16 //R5 = 10
		// mem[45] = 32'b1110_01_0_0100_1_0000_0110_000000010100; //LDR R6 ,[R0],#20 //R6 = 41	
		// mem[46] = 32'b1110_01_0_0100_1_0000_0111_000000011000; //LDR R7 ,[R0],#24 //R7 = 8912
		// mem[47] = 32'b1110_00_1_1101_0_0000_1000_000000000000; //MOV R8 ,#0 //R8 = 0
		// mem[48] = 32'b1110_00_1_1101_0_0000_1001_000000000000; //MOV R9 ,#0 //R9 = 0
		// mem[49] = 32'b1110_00_1_1101_0_0000_1010_000000000000; //MOV R10 ,#0 //R10 = 0
		// mem[50] = 32'b1110_00_1_1101_0_0000_1011_000000000000; //MOV R11 ,#0 //R11 = 0
		// mem[51] = 32'b1110_00_1_1101_0_0000_1100_000000000000; //MOV R12 ,#0 //R12 = 0
		// mem[52] = 32'b1110_00_1_1101_0_0000_1101_000000000000; //MOV R13 ,#0 //R13 = 0
		// mem[53] = 32'b1110_00_1_1101_0_0000_1110_000000000000; //MOV R14 ,#0 //R14 = 0
		// mem[54] = 32'b1110_10_1_0_111111111111111111111111 ;   //B #-1
		mem[27] = 32'b1110_10_1_0_111111111111111111111111 ;   //B #-1
	end
	
	assign Inst = mem[AddrIn[17:2]];

endmodule
