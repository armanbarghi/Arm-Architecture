module IF_Stage(input clk, rst, freeze, Branch_taken,
                input [31:0] BranchAddr,
                output reg [31:0] PC, Inst);

endmodule